-- Part_2_IF_ID.vhd
-- Implements the IF and ID blocks of a Simple Pipelined Architecture.

-- Design Phase 3
-- Date: 4/25/2025
-- Authors: Matthew Collins & Lewis Bates
-- Emails: mcollins42@tntech.edu & lfbates42@tntech.edu

library IEEE;
use IEEE.std_logic_1164.all;
use work.type_def.all;

-- Entity declaration for Part_2_IF_ID: Top-level module for IF and ID stages of a pipelined processor
entity Part_2_IF_ID is
    port (

        clk            : in  std_logic; 							-- Clock signal for synchronous operations
        reset          : in  std_logic; 							-- Reset signal to initialize registers
        branch_address : in  std_logic_vector(31 downto 0); -- Branch address input from EX stage for PC update
        pc_select      : in  std_logic; 							-- PC select signal to choose between normal or branch address
        write_register : in  std_logic_vector(4 downto 0); 	-- Write register address from WB stage for register file update
        write_data     : in  std_logic_vector(31 downto 0); -- Write data from WB stage to be stored in register file
        reg_write      : in  std_logic;         				-- Register write enable signal from WB stage
        
        -- Outputs to EX stage via ID/EX pipeline register
        ID_EX_PC_plus_4     : out std_logic_vector(31 downto 0); -- PC+4 value for EX stage
        ID_EX_rd_read_data  : out std_logic_vector(31 downto 0); -- Register rd read data
        ID_EX_rt_read_data  : out std_logic_vector(31 downto 0); -- Register rt read data
        ID_EX_sign_extended : out std_logic_vector(31 downto 0); -- Sign-extended immediate
        ID_EX_write_register: out std_logic_vector(4 downto 0);  -- Destination register address
        ID_EX_RegDst        : out std_logic;                     -- Register destination control signal
        ID_EX_Branch        : out std_logic;                     -- Branch control signal
        ID_EX_RegWrite      : out std_logic;                     -- Register write control signal
        ID_EX_ALUSrc        : out std_logic;                     -- ALU source control signal
        ID_EX_MemRead       : out std_logic;                     -- Memory read control signal
        ID_EX_MemWrite      : out std_logic;                     -- Memory write control signal
        ID_EX_MemtoReg      : out std_logic;                     -- Memory-to-register control signal
        ID_EX_ALUOp         : out std_logic_vector(1 downto 0)   -- ALU operation control signal
    );
end Part_2_IF_ID;

architecture Behavioral of Part_2_IF_ID is
    -- Component declarations for submodules used in IF and ID stages

    -- Program Counter (PC) component to store and update the current address
    component PC is
        port (
            Clock  	: in  std_logic;                     -- Clock input
            Resetn 	: in  std_logic;                     -- Reset input
            D  		: in  std_logic_vector(31 downto 0); -- Input PC value
            Q 			: out std_logic_vector(31 downto 0)  -- Output PC value
        );
    end component;

    -- Instruction memory component (single-port RAM) for fetching instructions
    component memory_1 is
        port (
            address : in  std_logic_vector(7 downto 0);  -- Memory address (byte-addressable)
            clock   : in  std_logic;                     -- Clock input
            data    : in  std_logic_vector(31 downto 0); -- Data input (not used here)
            wren    : in  std_logic;                     -- Write enable (not used here)
            q       : out std_logic_vector(31 downto 0)  -- Instruction output
        );
    end component;

    -- Multiplexer component to select between PC+4 and branch address
    component ALU_Mux is
        port (
            Input0 : in  std_logic_vector(31 downto 0); -- First input (PC+4)
            Input1 : in  std_logic_vector(31 downto 0); -- Second input (branch address)
            Sel    : in  std_logic;                     -- Select signal
            Output : out std_logic_vector(31 downto 0)  -- Selected output
        );
    end component;

    -- Control unit component to generate control signals based on opcode
    component control_unit is
        port (
            opcode   : in  std_logic_vector(5 downto 0);  -- Instruction opcode
            RegDst   : out std_logic;                     -- Register destination signal
            Branch   : out std_logic;                     -- Branch signal
            RegWrite : out std_logic;                     -- Register write signal
            ALUSrc   : out std_logic;                     -- ALU source signal
            MemRead  : out std_logic;                     -- Memory read signal
            MemWrite : out std_logic;                     -- Memory write signal
            MemtoReg : out std_logic;                     -- Memory-to-register signal
            ALUOp    : out std_logic_vector(1 downto 0)   -- ALU operation signal
        );
    end component;

    -- Register file component to store and access 32 registers
    component register_file is
       	port(
				read_reg_1		: IN STD_LOGIC_VECTOR(4 DOWNTO 0);		-- Read Register 1 Selection
				read_reg_2		: IN STD_LOGIC_VECTOR(4 DOWNTO 0);		-- Read Register 2 Selection
				write_reg		: IN STD_LOGIC_VECTOR(4 DOWNTO 0);		-- Write Register Selection
				write_data		: IN STD_LOGIC_VECTOR(31 DOWNTO 0);		-- Data to write to register
				regwrite_bit	: IN STD_LOGIC;								-- Enable Write
				reset				: IN STD_LOGIC;
				clock				: IN STD_LOGIC;
				read_data_1		: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);	-- Data stored in Read Register 1
				read_data_2		: OUT STD_LOGIC_VECTOR(31 DOWNTO 0) 	-- Data stored in Read register 2
			);
    end component;

    -- Sign extension component to extend 16-bit immediate to 32 bits
    component SignExtend is
        port (
            input  : in  std_logic_vector(15 downto 0);  -- 16-bit immediate input
            output : out std_logic_vector(31 downto 0)   -- 32-bit sign-extended output
        );
    end component;
	 
	 component pc_adder IS
    PORT (
        A : IN  STD_LOGIC_VECTOR(31 DOWNTO 0);  -- 32-bit input from PC
        B : IN  STD_LOGIC_VECTOR(31 DOWNTO 0);  -- 32-bit constant input (4)
        F : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)   -- 32-bit output (A + B)
    );
	 end component pc_adder;

    -- Internal signals for Instruction Fetch (IF) stage
    signal pc_current    : std_logic_vector(31 downto 0); -- Current program counter value
    signal pc_plus_4     : std_logic_vector(31 downto 0); -- PC incremented by 4
    signal instruction   : std_logic_vector(31 downto 0); -- Fetched instruction from memory
    signal mux1_out      : std_logic_vector(31 downto 0); -- Output of PC selection mux

    -- Internal signals for IF/ID pipeline register
    signal IF_ID_instruction : std_logic_vector(31 downto 0); -- Instruction stored in IF/ID register
    signal IF_ID_PC_plus_4   : std_logic_vector(31 downto 0); -- PC+4 stored in IF/ID register

    -- Internal signals for Instruction Decode (ID) stage
    signal reg_dst, branch, reg_write_id, alu_src, mem_read, mem_write, mem_to_reg : std_logic; -- Control signals from control unit
    signal alu_op : std_logic_vector(1 downto 0);           -- ALU operation code from control unit
    signal read_data1, read_data2 : std_logic_vector(31 downto 0); -- Data read from register file
    signal sign_extended : std_logic_vector(31 downto 0);   -- Sign-extended immediate value
    signal write_register_selected : std_logic_vector(4 downto 0); -- Selected destination register (rt or rd)

    -- Internal signals for ID/EX pipeline register (outputs to EX stage)
    signal ID_EX_PC_plus_4_reg     : std_logic_vector(31 downto 0); -- PC+4 value for EX stage
    signal ID_EX_rt_read_data1      : std_logic_vector(31 downto 0); -- Register rt data for EX stage
    signal ID_EX_rd_read_data1      : std_logic_vector(31 downto 0); -- Register rd data for EX stage
    signal ID_EX_sign_extended_reg : std_logic_vector(31 downto 0); -- Sign-extended immediate for EX stage
    signal ID_EX_write_register_reg: std_logic_vector(4 downto 0);  -- Destination register for EX stage
    signal ID_EX_RegDst_reg        : std_logic;                     -- RegDst control signal for EX stage
    signal ID_EX_Branch_reg        : std_logic;                     -- Branch control signal for EX stage
    signal ID_EX_RegWrite_reg      : std_logic;                     -- RegWrite control signal for EX stage
    signal ID_EX_ALUSrc_reg        : std_logic;                     -- ALUSrc control signal for EX stage
    signal ID_EX_MemRead_reg       : std_logic;                     -- MemRead control signal for EX stage
    signal ID_EX_MemWrite_reg      : std_logic;                     -- MemWrite control signal for EX stage
    signal ID_EX_MemtoReg_reg      : std_logic;                     -- MemtoReg control signal for EX stage
    signal ID_EX_ALUOp_reg         : std_logic_vector(1 downto 0);  -- ALUOp control signal for EX stage

begin
    -- Instruction Fetch (IF) Stage
    PC_inst : PC port map(
        Clock   => clk,          -- Clock signal for synchronization
        Resetn  => reset,        -- Reset signal to clear PC
        D       => mux1_out,     -- Next PC value from multiplexer
        Q       => pc_current    -- Current PC value output
    );

    adder_inst : pc_adder port map(
        A       => pc_current,   -- Matches pc_adder entity
        B       => "00000000000000000000000000000100", -- Constant 4
        F       => pc_plus_4     -- Matches pc_adder entity
    );

    instr_mem_inst : memory_1 port map(
        address => pc_current(7 downto 0),	-- Use lower 8 bits of PC as address
        clock   => clk,								-- Clock signal for memory access
        data    => (others => '0'),				-- Data input (unused for fetch)
        wren    => '0',								-- Write enable set to 0 (read-only)
        q       => instruction					-- Output fetched instruction
    );

    mux1_inst : ALU_Mux port map(
        Input0 => pc_plus_4,						-- Normal next PC (PC + 4)
        Input1 => branch_address,				-- Branch target address from EX stage
        Sel    => pc_select,						-- Selection signal from EX stage
        Output => mux1_out							-- Selected next PC valuec
    );

    -- IF/ID Pipeline Register: Latches IF stage outputs for ID stage
    process(clk)
    begin
        if rising_edge(clk) then
            if reset = '1' then
                -- Reset IF/ID register contents on reset
                IF_ID_instruction <= (others => '0');
                IF_ID_PC_plus_4   <= (others => '0');
            else
                -- Latch instruction and PC+4 on clock edge
                IF_ID_instruction <= instruction;
                IF_ID_PC_plus_4   <= pc_plus_4;
            end if;
        end if;
    end process;

    -- Instruction Decode (ID) Stage: Decodes instruction and prepares operands

    -- Instantiate control unit to generate control signals based on opcode
    control_unit_inst : control_unit port map(
        opcode   => IF_ID_instruction(31 downto 26), -- Opcode from fetched instruction
        RegDst   => reg_dst,                         -- Register destination signal
        Branch   => branch,                          -- Branch signal
        RegWrite => reg_write_id,                    -- Register write signal
        ALUSrc   => alu_src,                         -- ALU source signal
        MemRead  => mem_read,                        -- Memory read signal
        MemWrite => mem_write,                       -- Memory write signal
        MemtoReg => mem_to_reg,                      -- Memory-to-register signal
        ALUOp    => alu_op                           -- ALU operation signal
    );



    -- Instantiate register file to read source registers and write from WB stage
    register_file_inst : register_file port map(
		  read_reg_1	=> IF_ID_instruction(25 downto 21),		-- rs (source register 1)
		  read_reg_2	=> IF_ID_instruction(20 downto 16),		-- rt (source register 2)
		  write_reg		=> write_register,             			-- Write register from WB stage
		  write_data	=> write_data,                		   -- Write data from WB stage
		  regwrite_bit => reg_write,							  	   -- Write enable from WB stage
		  reset			=> reset,					   			   -- Reset signal
		  clock			=> clk,                           	   -- Clock signal for synchronization
		  read_data_1	=> read_data1,                         -- Data from rs
		  read_data_2	=> read_data2                          -- Data from rt	  
    );

    -- Instantiate sign extension unit to extend 16-bit immediate to 32 bits
    sign_extend_inst : SignExtend port map(
        input  => IF_ID_instruction(15 downto 0), -- 16-bit immediate from instruction
        output => sign_extended                   -- 32-bit sign-extended output
    );

    -- ID/EX Pipeline Register: Latches ID stage outputs for EX stage
    process(clk)
    begin
        if rising_edge(clk) then
            if reset = '1' then
                -- Reset ID/EX register contents on reset
                ID_EX_PC_plus_4_reg      <= (others => '0');
                ID_EX_rd_read_data1      <= (others => '0');
                ID_EX_rt_read_data1      <= (others => '0');
                ID_EX_sign_extended_reg  <= (others => '0');
                ID_EX_write_register_reg <= (others => '0');
                ID_EX_RegDst_reg         <= '0';
                ID_EX_Branch_reg         <= '0';
                ID_EX_RegWrite_reg       <= '0';
                ID_EX_ALUSrc_reg         <= '0';
                ID_EX_MemRead_reg        <= '0';
                ID_EX_MemWrite_reg       <= '0';
                ID_EX_MemtoReg_reg       <= '0';
                ID_EX_ALUOp_reg          <= (others => '0');
            else
                -- Latch ID stage outputs on clock edge for EX stage
                ID_EX_PC_plus_4_reg      <= IF_ID_PC_plus_4;         -- PC+4 value
                ID_EX_rd_read_data1      <= read_data1;              -- rd data
                ID_EX_rt_read_data1      <= read_data2;              -- rt data
                ID_EX_sign_extended_reg  <= sign_extended;           -- Sign-extended immediate
                ID_EX_write_register_reg <= write_register_selected; -- Destination register
                ID_EX_RegDst_reg         <= reg_dst;                 -- RegDst signal
                ID_EX_Branch_reg         <= branch;                  -- Branch signal
                ID_EX_RegWrite_reg       <= reg_write_id;            -- RegWrite signal
                ID_EX_ALUSrc_reg         <= alu_src;                 -- ALUSrc signal
                ID_EX_MemRead_reg        <= mem_read;                -- MemRead signal
                ID_EX_MemWrite_reg       <= mem_write;               -- MemWrite signal
                ID_EX_MemtoReg_reg       <= mem_to_reg;              -- MemtoReg signal
                ID_EX_ALUOp_reg          <= alu_op;                  -- ALUOp signal
            end if;
        end if;
    end process;

    -- Connect ID/EX register outputs to entity output ports for EX stage
    ID_EX_PC_plus_4     <= ID_EX_PC_plus_4_reg;      -- PC+4 to EX stage
    ID_EX_rd_read_data  <= ID_EX_rd_read_data1;       -- rd data to EX stage
    ID_EX_rt_read_data	<= ID_EX_rt_read_data1;       -- rt data to EX stage
    ID_EX_sign_extended <= ID_EX_sign_extended_reg;  -- Sign-extended immediate to EX stage
    ID_EX_write_register<= ID_EX_write_register_reg; -- Destination register to EX stage
    ID_EX_RegDst        <= ID_EX_RegDst_reg;         -- RegDst signal to EX stage
    ID_EX_Branch        <= ID_EX_Branch_reg;         -- Branch signal to EX stage
    ID_EX_RegWrite      <= ID_EX_RegWrite_reg;       -- RegWrite signal to EX stage
    ID_EX_ALUSrc        <= ID_EX_ALUSrc_reg;         -- ALUSrc signal to EX stage
    ID_EX_MemRead       <= ID_EX_MemRead_reg;        -- MemRead signal to EX stage
    ID_EX_MemWrite      <= ID_EX_MemWrite_reg;       -- MemWrite signal to EX stage
    ID_EX_MemtoReg      <= ID_EX_MemtoReg_reg;       -- MemtoReg signal to EX stage
    ID_EX_ALUOp         <= ID_EX_ALUOp_reg;          -- ALUOp signal to EX stage

end Behavioral;